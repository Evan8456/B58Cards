module player(
	input 
	output reg [9:0] hand // The memory address of the hand
	);

	initial begin
		hand = 0;
	end
endmodule
